SystemVerilog