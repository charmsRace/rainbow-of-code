Bluespec